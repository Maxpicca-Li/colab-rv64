`ifdef DEF_CONFIG
`define DEF_CONFIG

`define XLEN            64
`define REG_NUM         32
`define FIFO_CNT        16
`define REG_BUS         63:0
`define RST_PC          0

`endif